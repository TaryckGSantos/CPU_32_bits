- Fazer um set on less than pra ULA



Repositório para usar de parâmetro: https://github.com/dugagjin/MIPS/tree/master
