- Fazer um set on less than pra ULA
- Pesquisar como fazer o registerFile da maneira certa
- 


Repositório para usar de parâmetro: https://github.com/dugagjin/MIPS/tree/master
