- Fazer um set on less than pra ULA
